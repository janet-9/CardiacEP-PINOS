-80                 # Vm
-                   # Lambda
-                   # delLambda
-                   # Tension
-                   # Ke
-                   # Nae
-                   # Cae
7.05374e-13         # Iion
-                   # tension_component
-                   # illum
AlievPanfilovDynamic
0.0679341           # V

